module and_gate (
input wire and_in1,and_in2,
output wire and_out
);

assign and_out=and_in1 & and_in2;
endmodule