module reg_file(
input [4:0] a1,a2,a3,
input [31:0] write_data,
input clk,reset ,write_enable,
output [31:0] read_data1,read_data2
);
integer i;
reg [31:0] regster [31:0];
always @(posedge clk ,negedge reset)
    begin 
        if (!reset)
            for(i=0 ;i<31;i=i+1) 
                regster[i]<=32'h00000000;
            else if (write_enable)
                regster[a3]<=write_data;
    end 

assign read_data1=regster[a1];
assign read_data2=regster[a2];
endmodule 